interface  intf  () ;

    bit                    CLK               ;
    bit                    RST               ;
    bit [3:0]              SEED              ;
    bit                    OUT               ;
    bit                    Valid             ;
    
endinterface
